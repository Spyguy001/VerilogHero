module Main();

endmodule 